`timescale 1ns/1ns
module testbench();

reg A,B,C,D,E;
wire  ALARM;

mysource s (A,B,C,D,E,ALARM);

initial begin
    $dumpfile("TimingDiagram.vcd");
    $dumpvars(0,ALARM, A,B,C,D,E);
    A <= 0; B<= 0;C<=0;D<=0;E<=0;
#10 A <= 0; B<= 0;C<=0;D<=0;E<=1;
#10 A <= 0; B<= 0;C<=0;D<=1;E<=0;
#10 A <= 0; B<= 0;C<=0;D<=1;E<=1;
#10 A <= 0; B<= 0;C<=1;D<=0;E<=0;
#10 A <= 0; B<= 0;C<=1;D<=0;E<=1;
#10 A <= 0; B<= 0;C<=1;D<=1;E<=0;
#10 A <= 0; B<= 0;C<=1;D<=1;E<=1;
#10 A <= 0; B<= 1;C<=0;D<=0;E<=0;
#10 A <= 0; B<= 1;C<=0;D<=0;E<=1;
#10 A <= 0; B<= 1;C<=0;D<=1;E<=0;
#10 A <= 0; B<= 1;C<=0;D<=1;E<=1;
#10 A <= 0; B<= 1;C<=1;D<=0;E<=0;
#10 A <= 0; B<= 1;C<=1;D<=0;E<=1;
#10 A <= 0; B<= 1;C<=1;D<=1;E<=0;
#10 A <= 0; B<= 1;C<=1;D<=1;E<=1;
#10 A <= 1; B<= 0;C<=0;D<=0;E<=0;
#10 A <= 1; B<= 0;C<=0;D<=0;E<=1;
#10 A <= 1; B<= 0;C<=0;D<=1;E<=0;
#10 A <= 1; B<= 0;C<=0;D<=1;E<=1;
#10 A <= 1; B<= 0;C<=1;D<=0;E<=0;
#10 A <= 1; B<= 0;C<=1;D<=0;E<=1;
#10 A <= 1; B<= 0;C<=1;D<=1;E<=0;
#10 A <= 1; B<= 0;C<=1;D<=1;E<=1;
#10 A <= 1; B<= 1;C<=0;D<=0;E<=0;
#10 A <= 1; B<= 1;C<=0;D<=0;E<=1;
#10 A <= 1; B<= 1;C<=0;D<=1;E<=0;
#10 A <= 1; B<= 1;C<=0;D<=1;E<=1;
#10 A <= 1; B<= 1;C<=1;D<=0;E<=0;
#10 A <= 1; B<= 1;C<=1;D<=0;E<=1;
#10 A <= 1; B<= 1;C<=1;D<=1;E<=0;
#10 A <= 1; B<= 1;C<=1;D<=1;E<=1;
#10;

end

endmodule